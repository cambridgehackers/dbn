// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;
import Connectable::*;

// portz libraries
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import PortalMemory::*;

// generated by tool
import FpMacIndicationProxy::*;
import FpMacRequestWrapper::*;

// defined by user
import RbmTypes::*;
import FpMacTb::*;

module [Module] mkPortalTop(StdPortalTop#(addrWidth))
   provisos (Add#(a__, addrWidth, 40),
	     Add#(a__, b__, 40),
	     Add#(addrWidth, c__, 52),
	     Add#(addrWidth, d__, 64),
	     Add#(e__, f__, 40),
	     Add#(f__, 12, b__),
	     Add#(b__, g__, 44)
	     );

   FpMacIndicationProxy ind <- mkFpMacIndicationProxy(FpMacIndicationPortal);
   FpMacRequest req <- mkFpMacRequest(ind.ifc);
   FpMacRequestWrapper reqW <- mkFpMacRequestWrapper(FpMacRequestPortal,req);


   Vector#(2,StdPortal) portals;
   portals[0] = ind.portalIfc;
   portals[1] = reqW.portalIfc; 
   
   StdDirectory dir <- mkStdDirectory(portals);
   
   // when constructing ctrl and interrupt muxes, directories must be the first argument
   let ctrl_mux <- mkSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = nil;

endmodule : mkPortalTop
