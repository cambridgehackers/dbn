// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;
import Connectable::*;

// portz libraries
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import PortalMemory::*;
import MemServer::*;
import PortalMemory::*;
import Dma::*;
import DmaUtils::*;
import RbmTypes::*;

// generated by tool
import RbmRequestWrapper::*;
import MmRequestWrapper::*;
import SigmoidRequestWrapper::*;
import TimerRequestWrapper::*;
import DmaConfigWrapper::*;
import RbmIndicationProxy::*;
import MmIndicationProxy::*;
import SigmoidIndicationProxy::*;
import TimerIndicationProxy::*;
import DmaIndicationProxy::*;

// defined by user
import Rbm::*;

module [Module] mkPortalTop(PortalTop#(addrWidth,TMul#(32,N),Empty,1))
   provisos (Add#(a__, addrWidth, 40),
	     Add#(a__, b__, 40),
	     Add#(addrWidth, c__, 52),
	     Add#(addrWidth, d__, 64),
	     Add#(e__, f__, 40),
	     Add#(f__, 12, b__),
	     Add#(b__, g__, 44)
	     );

   DmaIndicationProxy dmaIndicationProxy <- mkDmaIndicationProxy(DmaIndicationPortal);

   RbmIndicationProxy rbmIndicationProxy <- mkRbmIndicationProxy(RbmIndicationPortal);
   MmIndicationProxy   mmIndicationProxy <- mkMmIndicationProxy(MmIndicationPortal);
   SigmoidIndicationProxy   sigmoidIndicationProxy <- mkSigmoidIndicationProxy(SigmoidIndicationPortal);
   TimerIndicationProxy timerIndicationProxy <- mkTimerIndicationProxy(TimerIndicationPortal);
   Rbm#(N) rbm <- mkRbm(rbmIndicationProxy.ifc, mmIndicationProxy.ifc, sigmoidIndicationProxy.ifc, timerIndicationProxy.ifc);
   RbmRequestWrapper rbmRequestWrapper <- mkRbmRequestWrapper(RbmRequestPortal,rbm.rbmRequest);
   MmRequestWrapper   mmRequestWrapper <- mkMmRequestWrapper(MmRequestPortal,rbm.mmRequest);
   SigmoidRequestWrapper   sigmoidRequestWrapper <- mkSigmoidRequestWrapper(SigmoidRequestPortal,rbm.sigmoidRequest);
   TimerRequestWrapper timerRequestWrapper <- mkTimerRequestWrapper(TimerRequestPortal,rbm.timerRequest);

   let readClients = rbm.readClients;
   Bool buffered = True;
   if (buffered) begin
      function Module#(DmaReadBuffer#(TMul#(N,32), 16)) mkBuffer(a x);
	 return mkDmaReadBuffer();
      endfunction
      let buffers <- mapM(mkBuffer, rbm.readClients);

      function Module#(Empty) connect(Tuple2#(DmaReadBuffer#(dsz, burstlen), ObjectReadClient#(dsz)) tpl);
	 return mkConnection(tpl_2(tpl), tpl_1(tpl).dmaServer);
      endfunction
      let connections <- mapM(connect, zip(buffers, rbm.readClients));

      function ObjectReadClient#(dsz) dmaClient(DmaReadBuffer#(dsz, burstlen) b);
	 return b.dmaClient;
      endfunction
      readClients = map(dmaClient, buffers);
   end
   else begin
      readClients = rbm.readClients;
   end

   let writeClients = rbm.writeClients;
   if (buffered) begin
      function Module#(DmaWriteBuffer#(TMul#(N,32), 16)) mkBuffer(a x);
	 return mkDmaWriteBuffer();
      endfunction
      let buffers <- mapM(mkBuffer, rbm.writeClients);

      function Module#(Empty) connect(Tuple2#(DmaWriteBuffer#(dsz, burstlen), ObjectWriteClient#(dsz)) tpl);
	 return mkConnection(tpl_2(tpl), tpl_1(tpl).dmaServer);
      endfunction
      let connections <- mapM(connect, zip(buffers, rbm.writeClients));

      function ObjectWriteClient#(dsz) dmaClient(DmaWriteBuffer#(dsz, burstlen) b);
	 return b.dmaClient;
      endfunction
      writeClients = map(dmaClient, buffers);
   end
   else begin
      writeClients = rbm.writeClients;
   end

   MemServer#(addrWidth, TMul#(32,N), 1) dma <- mkMemServer(dmaIndicationProxy.ifc, readClients, writeClients);

   DmaConfigWrapper dmaConfigWrapper <- mkDmaConfigWrapper(DmaConfigPortal,dma.request);

   Vector#(4,StdPortal) portals;
   portals[0] = rbmRequestWrapper.portalIfc;
   portals[1] = rbmIndicationProxy.portalIfc; 
   portals[2] = dmaConfigWrapper.portalIfc;
   portals[3] = dmaIndicationProxy.portalIfc; 
   
   StdDirectory dir <- mkStdDirectory(portals);
   
   // when constructing ctrl and interrupt muxes, directories must be the first argument
   let ctrl_mux <- mkSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;

endmodule : mkPortalTop
